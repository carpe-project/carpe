-- -*- vhdl -*-
-------------------------------------------------------------------------------
-- Copyright (c) 2012, The CARPE Project, All rights reserved.               --
-- See the AUTHORS file for individual contributors.                         --
--                                                                           --
-- Copyright and related rights are licensed under the Solderpad             --
-- Hardware License, Version 0.51 (the "License"); you may not use this      --
-- file except in compliance with the License. You may obtain a copy of      --
-- the License at http://solderpad.org/licenses/SHL-0.51.                    --
--                                                                           --
-- Unless required by applicable law or agreed to in writing, software,      --
-- hardware and materials distributed under this License is distributed      --
-- on an "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND,        --
-- either express or implied. See the License for the specific language      --
-- governing permissions and limitations under the License.                  --
-------------------------------------------------------------------------------


-- LRU Cache Replacement Algorithm

library ieee;
use ieee.std_logic_1164.all;

library util;
use util.numeric_pkg.all;

entity cache_replace_lru is

  generic (
    log2_assoc : natural := 1;
    index_bits : natural := 1
    );

  port (
    clk : in std_ulogic;
    rstn : in std_ulogic;

    re : in std_ulogic;
    rindex : in std_ulogic_vector(index_bits-1 downto 0);
    rway   : out std_ulogic_vector(2**log2_assoc-1 downto 0);
    rstate : out std_ulogic_vector((2**log2_assoc-1)*log2_assoc-1 downto 0);

    we : in std_ulogic;
    windex : in std_ulogic_vector(index_bits-1 downto 0);
    wway   : in std_ulogic_vector(2**log2_assoc-1 downto 0);
    wstate : in std_ulogic_vector((2**log2_assoc-1)*log2_assoc-1 downto 0)

    );
  
end;
